package tests_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import axi_if_pkg::*;
    import axi_env_pkg::*;

    `include "src/test_top.svh"
endpackage