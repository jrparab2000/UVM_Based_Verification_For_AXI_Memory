package axi_pkg_hdl;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    `include "src/axi_typedef.svh"
endpackage