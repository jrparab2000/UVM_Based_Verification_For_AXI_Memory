import uvm_pkg::*;
`include "uvm_macros.svh"
import tests_pkg::*;

module hvl_top ();
    initial begin
        run_test();
    end
endmodule