package tests_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import axi_if_pkg::*;
    import axi_env_pkg::*;
    import axi_sequences_pkg::*;
    `include "src/test_top.svh"
    `include "src/direct_test_seq_wr.svh"
endpackage